module test_module0 #(
	parameter      GROUP_NUM                      = 2       ,
	parameter      DW                             = 32      ,
	parameter      AW                             = 32      ,
	parameter      SW                             = 4       ,
	parameter      LW                             = 4       ,
	parameter      IDW                            = 6       ,
	parameter      AWUW                           = 16      ,
	parameter      ARUW                           = 16      ,
	parameter      RUW                            = 8       ,
	parameter      WUW                            = 4       ,
	parameter      BUW                            = 4       ,
	parameter      AW_TMO                         = 2       ,
	parameter      AR_TMO                         = 2       ,
	parameter      R_TMO                          = 2       ,
	parameter      W_TMO                          = 2       ,
	parameter      B_TMO                          = 2       ,
	localparam     DFX_AC                         = 1       ,
	localparam     RS_LTW                         = 1       ,
	localparam     RS_QOS_W                       = 4       ,
	parameter      MST_SLV                        = 0       ,
	parameter      CLAMP_SYNC                     = 0       ,
	parameter      CLAMP_ENABLE                   = 0       ,
	parameter      AWVLD_CLEN_TRANS_CYCLE_SRC     = 0       ,
	parameter      AWVLD_CLEN_TRANS_DELAY         = 0       ,
	parameter      AWVLD_CLEN_TRANS_CYCLE         = 1       ,
	parameter      AWVLD_CLEN_TRANS_RANDOM        = 1       ,
	parameter      AWVLD_CLEN_SYNC_RANDOM         = 1       ,
	parameter      ARVLD_CLEN_TRANS_CYCLE_SRC     = 0       ,
	parameter      ARVLD_CLEN_TRANS_DELAY         = 0       ,
	parameter      ARVLD_CLEN_TRANS_CYCLE         = 1       ,
	parameter      ARVLD_CLEN_TRANS_RANDOM        = 1       ,
	parameter      ARVLD_CLEN_SYNC_RANDOM         = 1       ,
	parameter      WVLD_CLEN_TRANS_CYCLE_SRC      = 0       ,
	parameter      WVLD_CLEN_TRANS_DELAY          = 0       ,
	parameter      WVLD_CLEN_TRANS_CYCLE          = 1       ,
	parameter      WVLD_CLEN_TRANS_RANDOM         = 1       ,
	parameter      WVLD_CLEN_SYNC_RANDOM          = 1       ,
	parameter      BVLD_CLEN_TRANS_CYCLE_SRC      = 0       ,
	parameter      BVLD_CLEN_TRANS_DELAY          = 0       ,
	parameter      BVLD_CLEN_TRANS_CYCLE          = 1       ,
	parameter      BVLD_CLEN_TRANS_RANDOM         = 1       ,
	parameter      BVLD_CLEN_SYNC_RANDOM          = 1       ,
	parameter      RVLD_CLEN_TRANS_CYCLE_SRC      = 0       ,
	parameter      RVLD_CLEN_TRANS_DELAY          = 0       ,
	parameter      RVLD_CLEN_TRANS_CYCLE          = 1       ,
	parameter      RVLD_CLEN_TRANS_RANDOM         = 1       ,
	parameter RVLD_CLEN_SYNC_RANDOM          = 1        
)(
input                                 aclk                     ,
input                                 aresetn                  ,
output  reg  [3:0]                    test_sig0_0              ,
output  reg  [3:0]                    test_sig0_1              ,
output  reg  [3:0]                    test_sig0_2              ,
output  reg  [3:0]                    test_sig0_3              ,
input        [EDF_MST_IDW-1:0]        mst_0_axi_awid           ,
input        [EDF_MST_AW-1:0]         mst_0_axi_awaddr         ,
input        [EDF_MST_LW-1:0]         mst_0_axi_awlen          ,
input        [2:0]                    mst_0_axi_awsize         ,
input        [1:0]                    mst_0_axi_awburst        ,
input                                 mst_0_axi_awlock         ,
input        [3:0]                    mst_0_axi_awcache        ,
input        [2:0]                    mst_0_axi_awprot         ,
input                                 mst_0_axi_awvalid        ,
output                                mst_0_axi_awready        ,
input        [EDF_MST_AWUW-1:0]       mst_0_axi_awuser         ,
input        [3:0]                    mst_0_axi_awqos          ,
input        [EDF_MST_IDW-1:0]        mst_0_axi_arid           ,
input        [EDF_MST_AW-1:0]         mst_0_axi_araddr         ,
input        [EDF_MST_LW-1:0]         mst_0_axi_arlen          ,
input        [2:0]                    mst_0_axi_arsize         ,
input        [1:0]                    mst_0_axi_arburst        ,
input                                 mst_0_axi_arlock         ,
input        [3:0]                    mst_0_axi_arcache        ,
input        [2:0]                    mst_0_axi_arprot         ,
input                                 mst_0_axi_arvalid        ,
output                                mst_0_axi_arready        ,
input        [EDF_MST_ARUW-1:0]       mst_0_axi_aruser         ,
input        [3:0]                    mst_0_axi_arqos          ,
input        [EDF_MST_DW-1:0]         mst_0_axi_wdata          ,
input        [EDF_MST_SW-1:0]         mst_0_axi_wstrb          ,
input                                 mst_0_axi_wlast          ,
input                                 mst_0_axi_wvalid         ,
output                                mst_0_axi_wready         ,
input        [EDF_MST_WUW-1:0]        mst_0_axi_wuser          ,
output       [EDF_MST_IDW-1:0]        mst_0_axi_bid            ,
output       [1:0]                    mst_0_axi_bresp          ,
output                                mst_0_axi_bvalid         ,
input                                 mst_0_axi_bready         ,
output       [EDF_MST_BUW-1:0]        mst_0_axi_buser          ,
output       [EDF_MST_IDW-1:0]        mst_0_axi_rid            ,
output       [EDF_MST_DW-1:0]         mst_0_axi_rdata          ,
output       [1:0]                    mst_0_axi_rresp          ,
output                                mst_0_axi_rlast          ,
output                                mst_0_axi_rvalid         ,
input                                 mst_0_axi_rready         ,
output       [EDF_MST_RUW-1:0]        mst_0_axi_ruser          ,
output       [EDF_MST_IDW-1:0]        slv_0_axi_awid           ,
output       [EDF_MST_AW-1:0]         slv_0_axi_awaddr         ,
output       [EDF_MST_LW-1:0]         slv_0_axi_awlen          ,
output       [2:0]                    slv_0_axi_awsize         ,
output       [1:0]                    slv_0_axi_awburst        ,
output                                slv_0_axi_awlock         ,
output       [3:0]                    slv_0_axi_awcache        ,
output       [2:0]                    slv_0_axi_awprot         ,
output                                slv_0_axi_awvalid        ,
input                                 slv_0_axi_awready        ,
output       [EDF_MST_AWUW-1:0]       slv_0_axi_awuser         ,
output       [3:0]                    slv_0_axi_awqos          ,
output       [EDF_MST_IDW-1:0]        slv_0_axi_arid           ,
output       [EDF_MST_AW-1:0]         slv_0_axi_araddr         ,
output       [EDF_MST_LW-1:0]         slv_0_axi_arlen          ,
output       [2:0]                    slv_0_axi_arsize         ,
output       [1:0]                    slv_0_axi_arburst        ,
output                                slv_0_axi_arlock         ,
output       [3:0]                    slv_0_axi_arcache        ,
output       [2:0]                    slv_0_axi_arprot         ,
output                                slv_0_axi_arvalid        ,
input                                 slv_0_axi_arready        ,
output       [EDF_MST_ARUW-1:0]       slv_0_axi_aruser         ,
output       [3:0]                    slv_0_axi_arqos          ,
output       [EDF_MST_DW-1:0]         slv_0_axi_wdata          ,
output       [EDF_MST_SW-1:0]         slv_0_axi_wstrb          ,
output                                slv_0_axi_wlast          ,
output                                slv_0_axi_wvalid         ,
input                                 slv_0_axi_wready         ,
output       [EDF_MST_WUW-1:0]        slv_0_axi_wuser          ,
input        [EDF_MST_IDW-1:0]        slv_0_axi_bid            ,
input        [1:0]                    slv_0_axi_bresp          ,
input                                 slv_0_axi_bvalid         ,
output                                slv_0_axi_bready         ,
input        [EDF_MST_BUW-1:0]        slv_0_axi_buser          ,
input        [EDF_MST_IDW-1:0]        slv_0_axi_rid            ,
input        [EDF_MST_DW-1:0]         slv_0_axi_rdata          ,
input        [1:0]                    slv_0_axi_rresp          ,
input                                 slv_0_axi_rlast          ,
input                                 slv_0_axi_rvalid         ,
output                                slv_0_axi_rready         ,
input        [EDF_MST_RUW-1:0]        slv_0_axi_ruser          ,
input        [EDF_MST_IDW-1:0]        mst_1_axi_awid           ,
input        [EDF_MST_AW-1:0]         mst_1_axi_awaddr         ,
input        [EDF_MST_LW-1:0]         mst_1_axi_awlen          ,
input        [2:0]                    mst_1_axi_awsize         ,
input        [1:0]                    mst_1_axi_awburst        ,
input                                 mst_1_axi_awlock         ,
input        [3:0]                    mst_1_axi_awcache        ,
input        [2:0]                    mst_1_axi_awprot         ,
input                                 mst_1_axi_awvalid        ,
output                                mst_1_axi_awready        ,
input        [EDF_MST_AWUW-1:0]       mst_1_axi_awuser         ,
input        [3:0]                    mst_1_axi_awqos          ,
input        [EDF_MST_IDW-1:0]        mst_1_axi_arid           ,
input        [EDF_MST_AW-1:0]         mst_1_axi_araddr         ,
input        [EDF_MST_LW-1:0]         mst_1_axi_arlen          ,
input        [2:0]                    mst_1_axi_arsize         ,
input        [1:0]                    mst_1_axi_arburst        ,
input                                 mst_1_axi_arlock         ,
input        [3:0]                    mst_1_axi_arcache        ,
input        [2:0]                    mst_1_axi_arprot         ,
input                                 mst_1_axi_arvalid        ,
output                                mst_1_axi_arready        ,
input        [EDF_MST_ARUW-1:0]       mst_1_axi_aruser         ,
input        [3:0]                    mst_1_axi_arqos          ,
input        [EDF_MST_DW-1:0]         mst_1_axi_wdata          ,
input        [EDF_MST_SW-1:0]         mst_1_axi_wstrb          ,
input                                 mst_1_axi_wlast          ,
input                                 mst_1_axi_wvalid         ,
output                                mst_1_axi_wready         ,
input        [EDF_MST_WUW-1:0]        mst_1_axi_wuser          ,
output       [EDF_MST_IDW-1:0]        mst_1_axi_bid            ,
output       [1:0]                    mst_1_axi_bresp          ,
output                                mst_1_axi_bvalid         ,
input                                 mst_1_axi_bready         ,
output       [EDF_MST_BUW-1:0]        mst_1_axi_buser          ,
output       [EDF_MST_IDW-1:0]        mst_1_axi_rid            ,
output       [EDF_MST_DW-1:0]         mst_1_axi_rdata          ,
output       [1:0]                    mst_1_axi_rresp          ,
output                                mst_1_axi_rlast          ,
output                                mst_1_axi_rvalid         ,
input                                 mst_1_axi_rready         ,
output       [EDF_MST_RUW-1:0]        mst_1_axi_ruser          ,
output       [EDF_MST_IDW-1:0]        slv_1_axi_awid           ,
output       [EDF_MST_AW-1:0]         slv_1_axi_awaddr         ,
output       [EDF_MST_LW-1:0]         slv_1_axi_awlen          ,
output       [2:0]                    slv_1_axi_awsize         ,
output       [1:0]                    slv_1_axi_awburst        ,
output                                slv_1_axi_awlock         ,
output       [3:0]                    slv_1_axi_awcache        ,
output       [2:0]                    slv_1_axi_awprot         ,
output                                slv_1_axi_awvalid        ,
input                                 slv_1_axi_awready        ,
output       [EDF_MST_AWUW-1:0]       slv_1_axi_awuser         ,
output       [3:0]                    slv_1_axi_awqos          ,
output       [EDF_MST_IDW-1:0]        slv_1_axi_arid           ,
output       [EDF_MST_AW-1:0]         slv_1_axi_araddr         ,
output       [EDF_MST_LW-1:0]         slv_1_axi_arlen          ,
output       [2:0]                    slv_1_axi_arsize         ,
output       [1:0]                    slv_1_axi_arburst        ,
output                                slv_1_axi_arlock         ,
output       [3:0]                    slv_1_axi_arcache        ,
output       [2:0]                    slv_1_axi_arprot         ,
output                                slv_1_axi_arvalid        ,
input                                 slv_1_axi_arready        ,
output       [EDF_MST_ARUW-1:0]       slv_1_axi_aruser         ,
output       [3:0]                    slv_1_axi_arqos          ,
output       [EDF_MST_DW-1:0]         slv_1_axi_wdata          ,
output       [EDF_MST_SW-1:0]         slv_1_axi_wstrb          ,
output                                slv_1_axi_wlast          ,
output                                slv_1_axi_wvalid         ,
input                                 slv_1_axi_wready         ,
output       [EDF_MST_WUW-1:0]        slv_1_axi_wuser          ,
input        [EDF_MST_IDW-1:0]        slv_1_axi_bid            ,
input        [1:0]                    slv_1_axi_bresp          ,
input                                 slv_1_axi_bvalid         ,
output                                slv_1_axi_bready         ,
input        [EDF_MST_BUW-1:0]        slv_1_axi_buser          ,
input        [EDF_MST_IDW-1:0]        slv_1_axi_rid            ,
input        [EDF_MST_DW-1:0]         slv_1_axi_rdata          ,
input        [1:0]                    slv_1_axi_rresp          ,
input                                 slv_1_axi_rlast          ,
input                                 slv_1_axi_rvalid         ,
output                                slv_1_axi_rready         ,
input        [EDF_MST_RUW-1:0]        slv_1_axi_ruser          ,
input        [EDF_MST_IDW-1:0]        mst_2_axi_awid           ,
input        [EDF_MST_AW-1:0]         mst_2_axi_awaddr         ,
input        [EDF_MST_LW-1:0]         mst_2_axi_awlen          ,
input        [2:0]                    mst_2_axi_awsize         ,
input        [1:0]                    mst_2_axi_awburst        ,
input                                 mst_2_axi_awlock         ,
input        [3:0]                    mst_2_axi_awcache        ,
input        [2:0]                    mst_2_axi_awprot         ,
input                                 mst_2_axi_awvalid        ,
output                                mst_2_axi_awready        ,
input        [EDF_MST_AWUW-1:0]       mst_2_axi_awuser         ,
input        [3:0]                    mst_2_axi_awqos          ,
input        [EDF_MST_IDW-1:0]        mst_2_axi_arid           ,
input        [EDF_MST_AW-1:0]         mst_2_axi_araddr         ,
input        [EDF_MST_LW-1:0]         mst_2_axi_arlen          ,
input        [2:0]                    mst_2_axi_arsize         ,
input        [1:0]                    mst_2_axi_arburst        ,
input                                 mst_2_axi_arlock         ,
input        [3:0]                    mst_2_axi_arcache        ,
input        [2:0]                    mst_2_axi_arprot         ,
input                                 mst_2_axi_arvalid        ,
output                                mst_2_axi_arready        ,
input        [EDF_MST_ARUW-1:0]       mst_2_axi_aruser         ,
input        [3:0]                    mst_2_axi_arqos          ,
input        [EDF_MST_DW-1:0]         mst_2_axi_wdata          ,
input        [EDF_MST_SW-1:0]         mst_2_axi_wstrb          ,
input                                 mst_2_axi_wlast          ,
input                                 mst_2_axi_wvalid         ,
output                                mst_2_axi_wready         ,
input        [EDF_MST_WUW-1:0]        mst_2_axi_wuser          ,
output       [EDF_MST_IDW-1:0]        mst_2_axi_bid            ,
output       [1:0]                    mst_2_axi_bresp          ,
output                                mst_2_axi_bvalid         ,
input                                 mst_2_axi_bready         ,
output       [EDF_MST_BUW-1:0]        mst_2_axi_buser          ,
output       [EDF_MST_IDW-1:0]        mst_2_axi_rid            ,
output       [EDF_MST_DW-1:0]         mst_2_axi_rdata          ,
output       [1:0]                    mst_2_axi_rresp          ,
output                                mst_2_axi_rlast          ,
output                                mst_2_axi_rvalid         ,
input                                 mst_2_axi_rready         ,
output       [EDF_MST_RUW-1:0]        mst_2_axi_ruser          ,
output       [EDF_MST_IDW-1:0]        slv_2_axi_awid           ,
output       [EDF_MST_AW-1:0]         slv_2_axi_awaddr         ,
output       [EDF_MST_LW-1:0]         slv_2_axi_awlen          ,
output       [2:0]                    slv_2_axi_awsize         ,
output       [1:0]                    slv_2_axi_awburst        ,
output                                slv_2_axi_awlock         ,
output       [3:0]                    slv_2_axi_awcache        ,
output       [2:0]                    slv_2_axi_awprot         ,
output                                slv_2_axi_awvalid        ,
input                                 slv_2_axi_awready        ,
output       [EDF_MST_AWUW-1:0]       slv_2_axi_awuser         ,
output       [3:0]                    slv_2_axi_awqos          ,
output       [EDF_MST_IDW-1:0]        slv_2_axi_arid           ,
output       [EDF_MST_AW-1:0]         slv_2_axi_araddr         ,
output       [EDF_MST_LW-1:0]         slv_2_axi_arlen          ,
output       [2:0]                    slv_2_axi_arsize         ,
output       [1:0]                    slv_2_axi_arburst        ,
output                                slv_2_axi_arlock         ,
output       [3:0]                    slv_2_axi_arcache        ,
output       [2:0]                    slv_2_axi_arprot         ,
output                                slv_2_axi_arvalid        ,
input                                 slv_2_axi_arready        ,
output       [EDF_MST_ARUW-1:0]       slv_2_axi_aruser         ,
output       [3:0]                    slv_2_axi_arqos          ,
output       [EDF_MST_DW-1:0]         slv_2_axi_wdata          ,
output       [EDF_MST_SW-1:0]         slv_2_axi_wstrb          ,
output                                slv_2_axi_wlast          ,
output                                slv_2_axi_wvalid         ,
input                                 slv_2_axi_wready         ,
output       [EDF_MST_WUW-1:0]        slv_2_axi_wuser          ,
input        [EDF_MST_IDW-1:0]        slv_2_axi_bid            ,
input        [1:0]                    slv_2_axi_bresp          ,
input                                 slv_2_axi_bvalid         ,
output                                slv_2_axi_bready         ,
input        [EDF_MST_BUW-1:0]        slv_2_axi_buser          ,
input        [EDF_MST_IDW-1:0]        slv_2_axi_rid            ,
input        [EDF_MST_DW-1:0]         slv_2_axi_rdata          ,
input        [1:0]                    slv_2_axi_rresp          ,
input                                 slv_2_axi_rlast          ,
input                                 slv_2_axi_rvalid         ,
output                                slv_2_axi_rready         ,
input        [EDF_MST_RUW-1:0]        slv_2_axi_ruser          ,
input        [EDF_MST_IDW-1:0]        mst_3_axi_awid           ,
input        [EDF_MST_AW-1:0]         mst_3_axi_awaddr         ,
input        [EDF_MST_LW-1:0]         mst_3_axi_awlen          ,
input        [2:0]                    mst_3_axi_awsize         ,
input        [1:0]                    mst_3_axi_awburst        ,
input                                 mst_3_axi_awlock         ,
input        [3:0]                    mst_3_axi_awcache        ,
input        [2:0]                    mst_3_axi_awprot         ,
input                                 mst_3_axi_awvalid        ,
output                                mst_3_axi_awready        ,
input        [EDF_MST_AWUW-1:0]       mst_3_axi_awuser         ,
input        [3:0]                    mst_3_axi_awqos          ,
input        [EDF_MST_IDW-1:0]        mst_3_axi_arid           ,
input        [EDF_MST_AW-1:0]         mst_3_axi_araddr         ,
input        [EDF_MST_LW-1:0]         mst_3_axi_arlen          ,
input        [2:0]                    mst_3_axi_arsize         ,
input        [1:0]                    mst_3_axi_arburst        ,
input                                 mst_3_axi_arlock         ,
input        [3:0]                    mst_3_axi_arcache        ,
input        [2:0]                    mst_3_axi_arprot         ,
input                                 mst_3_axi_arvalid        ,
output                                mst_3_axi_arready        ,
input        [EDF_MST_ARUW-1:0]       mst_3_axi_aruser         ,
input        [3:0]                    mst_3_axi_arqos          ,
input        [EDF_MST_DW-1:0]         mst_3_axi_wdata          ,
input        [EDF_MST_SW-1:0]         mst_3_axi_wstrb          ,
input                                 mst_3_axi_wlast          ,
input                                 mst_3_axi_wvalid         ,
output                                mst_3_axi_wready         ,
input        [EDF_MST_WUW-1:0]        mst_3_axi_wuser          ,
output       [EDF_MST_IDW-1:0]        mst_3_axi_bid            ,
output       [1:0]                    mst_3_axi_bresp          ,
output                                mst_3_axi_bvalid         ,
input                                 mst_3_axi_bready         ,
output       [EDF_MST_BUW-1:0]        mst_3_axi_buser          ,
output       [EDF_MST_IDW-1:0]        mst_3_axi_rid            ,
output       [EDF_MST_DW-1:0]         mst_3_axi_rdata          ,
output       [1:0]                    mst_3_axi_rresp          ,
output                                mst_3_axi_rlast          ,
output                                mst_3_axi_rvalid         ,
input                                 mst_3_axi_rready         ,
output       [EDF_MST_RUW-1:0]        mst_3_axi_ruser          ,
output       [EDF_MST_IDW-1:0]        slv_3_axi_awid           ,
output       [EDF_MST_AW-1:0]         slv_3_axi_awaddr         ,
output       [EDF_MST_LW-1:0]         slv_3_axi_awlen          ,
output       [2:0]                    slv_3_axi_awsize         ,
output       [1:0]                    slv_3_axi_awburst        ,
output                                slv_3_axi_awlock         ,
output       [3:0]                    slv_3_axi_awcache        ,
output       [2:0]                    slv_3_axi_awprot         ,
output                                slv_3_axi_awvalid        ,
input                                 slv_3_axi_awready        ,
output       [EDF_MST_AWUW-1:0]       slv_3_axi_awuser         ,
output       [3:0]                    slv_3_axi_awqos          ,
output       [EDF_MST_IDW-1:0]        slv_3_axi_arid           ,
output       [EDF_MST_AW-1:0]         slv_3_axi_araddr         ,
output       [EDF_MST_LW-1:0]         slv_3_axi_arlen          ,
output       [2:0]                    slv_3_axi_arsize         ,
output       [1:0]                    slv_3_axi_arburst        ,
output                                slv_3_axi_arlock         ,
output       [3:0]                    slv_3_axi_arcache        ,
output       [2:0]                    slv_3_axi_arprot         ,
output                                slv_3_axi_arvalid        ,
input                                 slv_3_axi_arready        ,
output       [EDF_MST_ARUW-1:0]       slv_3_axi_aruser         ,
output       [3:0]                    slv_3_axi_arqos          ,
output       [EDF_MST_DW-1:0]         slv_3_axi_wdata          ,
output       [EDF_MST_SW-1:0]         slv_3_axi_wstrb          ,
output                                slv_3_axi_wlast          ,
output                                slv_3_axi_wvalid         ,
input                                 slv_3_axi_wready         ,
output       [EDF_MST_WUW-1:0]        slv_3_axi_wuser          ,
input        [EDF_MST_IDW-1:0]        slv_3_axi_bid            ,
input        [1:0]                    slv_3_axi_bresp          ,
input                                 slv_3_axi_bvalid         ,
output                                slv_3_axi_bready         ,
input        [EDF_MST_BUW-1:0]        slv_3_axi_buser          ,
input        [EDF_MST_IDW-1:0]        slv_3_axi_rid            ,
input        [EDF_MST_DW-1:0]         slv_3_axi_rdata          ,
input        [1:0]                    slv_3_axi_rresp          ,
input                                 slv_3_axi_rlast          ,
input                                 slv_3_axi_rvalid         ,
output                                slv_3_axi_rready         ,
input        [EDF_MST_RUW-1:0]        slv_3_axi_ruser          
);
endmodule
